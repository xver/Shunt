`define MY_HOST "localhost"
`define MY_PORT  3450
`define V_SIZE   5
`define STRING_MESSAGE "server function int string_loopback_test(int socket_id)\0"
`define STRING_MESSAGE1 "SERVER FUNCTION INT STRING_LOOPBACK_TEST(INT SOCKET_ID)\0" 

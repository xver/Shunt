/*
 =========================================================
 File        : shunt_vcs_dpi.h
 Version     : 1.0.1
 Copyright (c) 2016-2017 IC Verimeter. All rights reserved.
 Licensed under the MIT License.
 See LICENSE file in the project root for full license information.
 Description : shunt vcs integration

 Not supported DPI functions defines:
 Version 1.0.1 : VCS

 System Verilog target initiator handshake (TCP/IP SystemVerilog SHUNT)
 ******************************************************
*/

`define NO_SHUNT_DPI_SEND_BITN
`define NO_SHUNT_DPI_RECV_BITN
`define NO_SHUNT_DPI_HS_SEND_BITN
`define NO_SHUNT_DPI_HS_RECV_BITN
`define NO_SHUNT_DPI_HS_SEND_REGN
`define NO_SHUNT_DPI_HS_SEND_LOGICN
`define NO_SHUNT_DPI_HS_RECV_REGN
`define NO_SHUNT_DPI_HS_RECV_LOGICN
`define NO_SHUNT_DPI_SEND_TIME
`define NO_SHUNT_DPI_RECV_TIME

`endif //  `ifndef SHUNT_VCS_DPI_H




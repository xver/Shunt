`define MY_HOST "localhost"
`define MY_PORT  3450


`define MY_HOST "localhost"
`define MY_PORT  3450
`define V_SIZE   5
 

